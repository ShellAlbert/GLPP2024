module ZCfgOV5640ByFPGA(
	input iClk,
	input iRST_N,
	input iStartPulse,
	output oDonePulse,
	output oI2C_SCL,
	inout ioI2C_SDA
);
endmodule
