module ZClkDivider4SCCB(
	input iClk,
	input iRst_N,
	input iEn,
	output oClk
);
endmodule