module ZCfgM3256LByFPGA(
	input iClk,
	input iRst_N,
	input iEn,
	output oCfgDone,
	output oUART_Txd,
	input iUART_Rxd
);

endmodule
