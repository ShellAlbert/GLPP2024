module ZCfgOV5640BySTM32(
	input iClk,
	input iRST_N,
	input iStartPulse,
	output oDonePulse,
	output oI2C_SCL,
	inout ioI2C_SDA
);
endmodule
